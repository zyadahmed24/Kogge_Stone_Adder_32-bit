
#******
# Preview export LEF
#
#	 Preview sub-version 5.10.41.500.3.38
#
# TECH LIB NAME: tsmc18
# TECH FILE NAME: techfile.cds
#******

VERSION 5.4 ;

NAMESCASESENSITIVE ON ;

DIVIDERCHAR "|" ;
BUSBITCHARS "[]" ;

UNITS
    DATABASE MICRONS 100  ;
END UNITS

MACRO KG_TOP
    CLASS CORE ;
    FOREIGN KG_TOP 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 120 BY 120 ;
    SYMMETRY X Y ;
    PIN A[0]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  2 95.00 2.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[0]
    PIN A[1]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  4 95.00 4.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[1]
    PIN A[2]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  6 95.00 6.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[2]
    PIN A[3]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  8 95.00 8.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[3]
    PIN A[4]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  10 95.00 10.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[4]
    PIN A[5]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  12 95.00 12.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[5]
    PIN A[6]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  14 95.00 14.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[6]
    PIN A[7]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  16 95.00 16.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[7]
    PIN A[8]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  18 95.00 18.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[8]
    PIN A[9]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  20 95.00 20.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[9]
    PIN A[10]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  22 95.00 22.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[10]
    PIN A[11]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  24 95.00 24.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[11]
    PIN A[12]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  26 95.00 26.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[12]
    PIN A[13]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  28 95.00 28.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[13]
    PIN A[14]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  30 95.00 30.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[14]
    PIN A[15]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  32 95.00 32.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[15]
    PIN A[16]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  34 95.00 34.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[16]
    PIN A[17]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  36 95.00 36.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[17]
    PIN A[18]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  38 95.00 38.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[18]
    PIN A[19]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  40 95.00 40.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[19]
    PIN A[20]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  42 95.00 42.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[20]
    PIN A[21]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  44 95.00 44.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[21]
    PIN A[22]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  46 95.00 46.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[22]
    PIN A[23]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  48 95.00 48.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[23]
    PIN A[24]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  50 95.00 50.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[24]
    PIN A[25]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  52 95.00 52.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[25]
    PIN A[26]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  54 95.00 54.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[26]
    PIN A[27]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  56 95.00 56.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[27]
    PIN A[28]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  58 95.00 58.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[28]
    PIN A[29]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  60 95.00 60.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[29]
    PIN A[30]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  62 95.00 62.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[30]
    PIN A[31]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  64 95.00 64.2 95.2 ;
        END
	AntennaGateArea 0.0 ;
    END A[31]
    PIN B[0]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 11 0.2 11.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[0]
    PIN B[1]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 13 0.2 13.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[1]
    PIN B[2]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 15 0.2 15.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[2]
    PIN B[3]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 17 0.2 17.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[3]
    PIN B[4]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 19 0.2 19.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[4]
    PIN B[5]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 21 0.2 21.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[5]
    PIN B[6]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 23 0.2 23.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[6]
    PIN B[7]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 25 0.2 25.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[7]
    PIN B[8]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 27 0.2 27.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[8]
    PIN B[9]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 29 0.2 29.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[9]
    PIN B[10]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 31 0.2 31.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[10]
    PIN B[11]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 33 0.2 33.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[11]
    PIN B[12]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 35 0.2 35.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[12]
    PIN B[13]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 37 0.2 37.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[13]
    PIN B[14]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 39 0.2 39.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[14]
    PIN B[15]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 41 0.2 41.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[15]
    PIN B[16]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 43 0.2 43.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[16]
    PIN B[17]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 45 0.2 45.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[17]
    PIN B[18]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 47 0.2 47.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[18]
    PIN B[19]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 49 0.2 49.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[19]
    PIN B[20]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 51 0.2 51.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[20]
    PIN B[21]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 53 0.2 53.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[21]
    PIN B[22]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 55 0.2 55.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[22]
    PIN B[23]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 57 0.2 57.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[23]
    PIN B[24]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 59 0.2 59.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[24]
    PIN B[25]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 61 0.2 61.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[25]
    PIN B[26]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 63 0.2 63.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[26]
    PIN B[27]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 65 0.2 65.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[27]
    PIN B[28]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 67 0.2 67.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[28]
    PIN B[29]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 69 0.2 69.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[29]
    PIN B[30]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 71 0.2 71.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[30]
    PIN B[31]
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 73 0.2 73.2 ;
        END
	AntennaGateArea 0.0 ;
    END B[31]
    PIN Cin
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 70 0.2 70.2 ;
        END
	AntennaGateArea 0.0 ;
    END Cin
    PIN clk
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 74 0.2 74.2 ;
        END
	AntennaGateArea 0.0 ;
    END clk
    PIN rst
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.00 78 0.2 78.2 ;
        END
	AntennaGateArea 0.0 ;
    END rst
    PIN S[0]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 2 95.2 2.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[0]
    PIN S[1]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 4 95.2 4.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[1]
    PIN S[2]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 6 95.2 6.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[2]
    PIN S[3]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 8 95.2 8.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[3]
    PIN S[4]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 10 95.2 10.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[4]
    PIN S[5]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 12 95.2 12.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[5]
    PIN S[6]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 14 95.2 14.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[6]
    PIN S[7]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 16 95.2 16.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[7]
    PIN S[8]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 18 95.2 18.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[8]
    PIN S[9]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 20 95.2 20.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[9]
    PIN S[10]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 22 95.2 22.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[10]
    PIN S[11]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 24 95.2 24.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[11]
    PIN S[12]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 26 95.2 26.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[12]
    PIN S[13]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 28 95.2 28.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[13]
    PIN S[14]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 30 95.2 30.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[14]
    PIN S[15]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 32 95.2 32.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[15]
    PIN S[16]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 34 95.2 34.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[16]
    PIN S[17]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 36 95.2 36.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[17]
    PIN S[18]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 38 95.2 38.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[18]
    PIN S[19]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 40 95.2 40.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[19]
    PIN S[20]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 42 95.2 42.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[20]
    PIN S[21]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 44 95.2 44.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[21]
    PIN S[22]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 46 95.2 46.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[22]
    PIN S[23]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 48 95.2 48.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[23]
    PIN S[24]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 50 95.2 50.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[24]
    PIN S[25]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 52 95.2 52.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[25]
    PIN S[26]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 54 95.2 54.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[26]
    PIN S[27]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 56 95.2 56.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[27]
    PIN S[28]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 58 95.2 58.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[28]
    PIN S[29]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 60 95.2 60.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[29]
    PIN S[30]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 62 95.2 62.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[30]
    PIN S[31]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 64 95.2 64.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[31]
    PIN S[32]
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  95.00 66 95.2 66.2 ;
        END
	AntennaGateArea 0.0 ;
    END S[32]
    END KG_TOP

END LIBRARY

