module dff_out #(parameter OUTPUT_WIDTH = 33) (
	input wire clk, rst,
	input wire [OUTPUT_WIDTH-1:0] S_D,
	
	output reg [OUTPUT_WIDTH-1:0] S_Q
);

always @(posedge clk or negedge rst) begin
	if(!rst) begin
		S_Q <= 'b0;
	end
	else begin
		S_Q <= S_D;
	end
end

endmodule
